// maoin_tb.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module maoin_tb (
	);

	wire    maoin_inst_clk_bfm_clk_clk;       // maoin_inst_clk_bfm:clk -> [maoin_inst:clk_clk, maoin_inst_reset_bfm:clk]
	wire    maoin_inst_reset_bfm_reset_reset; // maoin_inst_reset_bfm:reset -> maoin_inst:reset_reset_n

	maoin maoin_inst (
		.clk_clk       (maoin_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (maoin_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) maoin_inst_clk_bfm (
		.clk (maoin_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) maoin_inst_reset_bfm (
		.reset (maoin_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (maoin_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
