
module maoin (
	btn0_i_export,
	clk_clk,
	led0_o_export,
	reset_reset_n);	

	input		btn0_i_export;
	input		clk_clk;
	output	[7:0]	led0_o_export;
	input		reset_reset_n;
endmodule
